`timescale 1ns / 1ps

module top (
    (* dont_touch = "true" *)
    input  wire          clk100,
    output wire          serial_tx,
    input  wire          serial_rx,
    output wire          lpddr4_clk_p,
    output wire          lpddr4_clk_n,
    output wire          lpddr4_cke,
    output wire          lpddr4_odt,
    output wire          lpddr4_reset_n,
    output wire          lpddr4_cs,
    output wire    [5:0] lpddr4_ca,
    inout  wire   [15:0] lpddr4_dq,
    inout  wire    [1:0] lpddr4_dqs_p,
    inout  wire    [1:0] lpddr4_dqs_n,
    inout  wire    [1:0] lpddr4_dmi,
    output wire          user_led0,
    output wire          user_led1,
    output wire          user_led2,
    output wire          user_led3,
    output wire          user_led4,
    input  wire          user_btn0,
    input  wire          user_btn1
);

dram_phy phy_inst (
    .serial_tx(serial_tx),
    .serial_rx(serial_rx),
    .clk(clk100),
    .rst(~user_btn0),
    .clk_idelay(),
    .rst_idelay(),
    .clk_sys(),
    .rst_sys(),
    .clk_sys2x(),
    .rst_sys2x(),
    .clk_sys8x(),
    .rst_sys8x(),
    .ddram_ca(lpddr4_ca),
    .ddram_cs(lpddr4_cs),
    .ddram_dq(lpddr4_dq),
    .ddram_dqs_p(lpddr4_dqs_p),
    .ddram_dqs_n(lpddr4_dqs_n),
    .ddram_dmi(lpddr4_dmi),
    .ddram_clk_p(lpddr4_clk_p),
    .ddram_clk_n(lpddr4_clk_n),
    .ddram_cke(lpddr4_cke),
    .ddram_odt(lpddr4_odt),
    .ddram_reset_n(lpddr4_reset_n),
    .dfi_cke_p0(),
    .dfi_reset_n_p0(),
    .dfi_mode_2n_p0(),
    .dfi_alert_n_w0(),
    .dfi_address_p0(),
    .dfi_bank_p0(),
    .dfi_cas_n_p0(),
    .dfi_cs_n_p0(),
    .dfi_ras_n_p0(),
    .dfi_act_n_p0(),
    .dfi_odt_p0(),
    .dfi_we_n_p0(),
    .dfi_wrdata_p0(),
    .dfi_wrdata_en_p0(),
    .dfi_wrdata_mask_p0(),
    .dfi_rddata_en_p0(),
    .dfi_rddata_w0(),
    .dfi_rddata_valid_w0(),
    .dfi_cke_p1(),
    .dfi_reset_n_p1(),
    .dfi_mode_2n_p1(),
    .dfi_alert_n_w1(),
    .dfi_address_p1(),
    .dfi_bank_p1(),
    .dfi_cas_n_p1(),
    .dfi_cs_n_p1(),
    .dfi_ras_n_p1(),
    .dfi_act_n_p1(),
    .dfi_odt_p1(),
    .dfi_we_n_p1(),
    .dfi_wrdata_p1(),
    .dfi_wrdata_en_p1(),
    .dfi_wrdata_mask_p1(),
    .dfi_rddata_en_p1(),
    .dfi_rddata_w1(),
    .dfi_rddata_valid_w1(),
    .dfi_cke_p2(),
    .dfi_reset_n_p2(),
    .dfi_mode_2n_p2(),
    .dfi_alert_n_w2(),
    .dfi_address_p2(),
    .dfi_bank_p2(),
    .dfi_cas_n_p2(),
    .dfi_cs_n_p2(),
    .dfi_ras_n_p2(),
    .dfi_act_n_p2(),
    .dfi_odt_p2(),
    .dfi_we_n_p2(),
    .dfi_wrdata_p2(),
    .dfi_wrdata_en_p2(),
    .dfi_wrdata_mask_p2(),
    .dfi_rddata_en_p2(),
    .dfi_rddata_w2(),
    .dfi_rddata_valid_w2(),
    .dfi_cke_p3(),
    .dfi_reset_n_p3(),
    .dfi_mode_2n_p3(),
    .dfi_alert_n_w3(),
    .dfi_address_p3(),
    .dfi_bank_p3(),
    .dfi_cas_n_p3(),
    .dfi_cs_n_p3(),
    .dfi_ras_n_p3(),
    .dfi_act_n_p3(),
    .dfi_odt_p3(),
    .dfi_we_n_p3(),
    .dfi_wrdata_p3(),
    .dfi_wrdata_en_p3(),
    .dfi_wrdata_mask_p3(),
    .dfi_rddata_en_p3(),
    .dfi_rddata_w3(),
    .dfi_rddata_valid_w3(),
    .dfi_cke_p4(),
    .dfi_reset_n_p4(),
    .dfi_mode_2n_p4(),
    .dfi_alert_n_w4(),
    .dfi_address_p4(),
    .dfi_bank_p4(),
    .dfi_cas_n_p4(),
    .dfi_cs_n_p4(),
    .dfi_ras_n_p4(),
    .dfi_act_n_p4(),
    .dfi_odt_p4(),
    .dfi_we_n_p4(),
    .dfi_wrdata_p4(),
    .dfi_wrdata_en_p4(),
    .dfi_wrdata_mask_p4(),
    .dfi_rddata_en_p4(),
    .dfi_rddata_w4(),
    .dfi_rddata_valid_w4(),
    .dfi_cke_p5(),
    .dfi_reset_n_p5(),
    .dfi_mode_2n_p5(),
    .dfi_alert_n_w5(),
    .dfi_address_p5(),
    .dfi_bank_p5(),
    .dfi_cas_n_p5(),
    .dfi_cs_n_p5(),
    .dfi_ras_n_p5(),
    .dfi_act_n_p5(),
    .dfi_odt_p5(),
    .dfi_we_n_p5(),
    .dfi_wrdata_p5(),
    .dfi_wrdata_en_p5(),
    .dfi_wrdata_mask_p5(),
    .dfi_rddata_en_p5(),
    .dfi_rddata_w5(),
    .dfi_rddata_valid_w5(),
    .dfi_cke_p6(),
    .dfi_reset_n_p6(),
    .dfi_mode_2n_p6(),
    .dfi_alert_n_w6(),
    .dfi_address_p6(),
    .dfi_bank_p6(),
    .dfi_cas_n_p6(),
    .dfi_cs_n_p6(),
    .dfi_ras_n_p6(),
    .dfi_act_n_p6(),
    .dfi_odt_p6(),
    .dfi_we_n_p6(),
    .dfi_wrdata_p6(),
    .dfi_wrdata_en_p6(),
    .dfi_wrdata_mask_p6(),
    .dfi_rddata_en_p6(),
    .dfi_rddata_w6(),
    .dfi_rddata_valid_w6(),
    .dfi_cke_p7(),
    .dfi_reset_n_p7(),
    .dfi_mode_2n_p7(),
    .dfi_alert_n_w7(),
    .dfi_address_p7(),
    .dfi_bank_p7(),
    .dfi_cas_n_p7(),
    .dfi_cs_n_p7(),
    .dfi_ras_n_p7(),
    .dfi_act_n_p7(),
    .dfi_odt_p7(),
    .dfi_we_n_p7(),
    .dfi_wrdata_p7(),
    .dfi_wrdata_en_p7(),
    .dfi_wrdata_mask_p7(),
    .dfi_rddata_en_p7(),
    .dfi_rddata_w7(),
    .dfi_rddata_valid_w7(),
    .dfi_init_start(~user_btn1),
    .dfi_init_complete(user_led0)
);

endmodule